`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: lab1
//////////////////////////////////////////////////////////////////////////////////


module lab1(
    input [15:0] a,
     output [15:0] b
    );
    
    assign b[0] = ~a[0];
    assign b[1] = a[1] & ~a[2];
    assign b[3] = a[2] & a[3];
    assign b[2] = b[1] | b[3];   
    assign b[15:4] = a[15:4];
    
endmodule
